// Ques. write verilog code for a module that has no input and a constant output at logic high

module top_module ( output one );
  assign one = 1'b1;
endmodule 
