module buffer_mod ( input in , output out);
  assign out = in;
endmodule
