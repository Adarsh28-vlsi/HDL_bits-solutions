// Ques. write a verilog code for a module with no inputs and one output constant at logic zero
module top_module( output zero );
  assign zero = 1'b0;
endmodule
